module Not16 (input [15:0] in,
              output [15:0] out);
   Not n0(.in(in[0]), .out(out[0]));
   Not n1(.in(in[1]), .out(out[1]));
   Not n2(.in(in[2]), .out(out[2]));
   Not n3(.in(in[3]), .out(out[3]));
   Not n4(.in(in[4]), .out(out[4]));
   Not n5(.in(in[5]), .out(out[5]));
   Not n6(.in(in[6]), .out(out[6]));
   Not n7(.in(in[7]), .out(out[7]));
   Not n8(.in(in[8]), .out(out[8]));
   Not n9(.in(in[9]), .out(out[9]));
   Not n10(.in(in[10]), .out(out[10]));
   Not n11(.in(in[11]), .out(out[11]));
   Not n12(.in(in[12]), .out(out[12]));
   Not n13(.in(in[13]), .out(out[13]));
   Not n14(.in(in[14]), .out(out[14]));
   Not n15(.in(in[15]), .out(out[15]));
endmodule
